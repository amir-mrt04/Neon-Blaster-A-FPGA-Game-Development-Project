library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.math_real.all;
entity VGA_Square is
  port ( CLK_24MHz		: in std_logic;
			RESET				: in std_logic;
			Btn          : in std_logic_vector(3 downto 0);  --use Key(0) to Btn
			end_game       : in bit;
			pause        : in bit;			
			score          : out integer;
			lose           : out bit;
			ColorOut			: out std_logic_vector(5 downto 0); 
			SQUAREWIDTH		: in std_logic_vector(7 downto 0);
			ScanlineX		: in std_logic_vector(10 downto 0);
			random : in integer range 0 to 24000000;
			ScanlineY		: in std_logic_vector(10 downto 0)
  );
end VGA_Square;

architecture Behavioral of VGA_Square is
  
  
  signal ColorOutput: std_logic_vector(5 downto 0);
  signal SquareX: std_logic_vector(9 downto 0):="1111111111";  
  signal SquareY: std_logic_vector(9 downto 0):="1111111111";  
  signal Prescaler: std_logic_vector(30 downto 0); 
  signal rockX: std_logic_vector(9 downto 0):="1111111111";
  signal rockY: std_logic_vector(9 downto 0):="1111111111";
  signal rocknum: integer range 0 to 9 :=3; 
  signal rockdam,savedam: integer range 0 to 9 :=3;
  signal rockflag,fast,losegame: bit := '0' ;
  signal speed: integer := 100000 ;
  signal shotX: std_logic_vector(9 downto 0):="1111111111";
  signal shotY: std_logic_vector(9 downto 0):="1111111111";
  signal shotsize: std_logic_vector(9 downto 0):="0000000111";
  signal score_signal: integer range 0 to 99 :=0;
  signal wall_color : std_logic_vector(5 downto 0);
  	type BITMAP is array (0 to 21, 0 to 21) of bit ;
	type BITMAP2 is array (0 to 6, 0 to 6) of bit ;
	type BITMAP3 is array (0 to 21, 0 to 65) of bit ;
	constant endWin: bitMap3 := (
	('0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1'),
	('1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1'),
	('1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1'),
	('1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0'),
	('0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0'),
	('0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0'),
	('0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0'),
	('0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0'),
	('0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0'),
	('0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0'),
	('0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0'),
	('0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0'),
	('0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0'),
	('0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0'),
	('0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0'),
	('0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0'),
	('0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0'),
	('0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0'),
	('0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'),
	('0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'),
	('0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'),	
	('0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0'));
	constant endlose : bitMap3 := (
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0'),
	('1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0'),
	('1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0'));


	constant shotmap : BITMAP2 :=(	('0','0','0','1','0','0','0'),
											('0','0','1','1','1','0','0'),
											('0','1','1','1','1','1','0'),
											('1','1','1','1','1','1','1'),
											('0','1','1','1','1','1','0'),
											('0','0','1','1','1','0','0'),
											('0','0','0','1','0','0','0'));
	signal rockmap :BITMAP ;
		constant rock1 : BITMAP :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
	('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));	
	constant rock2 : BITMAP :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));	
	constant rock3 : BITMAP :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));	
		constant rock4 : BITMAP :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
	constant rock5 : BITMAP :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));	
	constant rock6: BITMAP :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));	
		constant rock7 : BITMAP :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
	constant rock8 : BITMAP :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
constant tank : BITMAP :=(('0','0','0','0','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
constant wall : BITMAP := (('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0'),
('0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0'),
('0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0'),
('0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0'),
('0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0'),
('0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0'),
('0','1','1','0','0','0','0','0','0','1','0','0','1','0','0','0','0','0','0','1','1','0'),
('0','1','1','0','0','0','0','0','1','0','0','0','0','1','0','0','0','0','0','1','1','0'),
('0','1','1','0','0','0','0','1','0','0','0','0','0','0','1','0','0','0','0','1','1','0'),
('0','1','1','1','1','1','1','0','0','0','1','1','0','0','0','1','1','1','1','1','1','0'),
('0','1','1','1','1','1','1','0','0','0','1','1','0','0','0','1','1','1','1','1','1','0'),
('0','1','1','0','0','0','0','1','0','0','0','0','0','0','1','0','0','0','0','1','1','0'),
('0','1','1','0','0','0','0','0','1','0','0','0','0','1','0','0','0','0','0','1','1','0'),
('0','1','1','0','0','0','0','0','0','1','0','0','1','0','0','0','0','0','0','1','1','0'),
('0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0'),
('0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0'),
('0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0'),
('0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0'),
('0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0'),
('0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0'),
('0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0'));
		constant home : BITMAP :=(('0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0'),
('0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','1','0','0','0','0','0'),
('0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','1','0','0','0','0'),
('0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','0','0','0'),
('0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','0','0'),
('0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0'),
('0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','0','0','1','0'),
('0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','0','0','1','0'),
('0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','0','0','1','0'),
('0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','0'),
('0','1','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','1','0'),
('0','1','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','1','0'),
('0','1','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','1','0'),
('0','1','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','1','0'),
('0','1','0','1','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','1','0'),
('0','1','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','1','0'),
('0','1','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','1','0'),
('0','1','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','1','0'),
('0','1','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','1','0'),
('0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
begin

square: process(CLK_24MHz, RESET)
	variable flag_btn,flagR,flagL : bit := '0';
	variable lock_key: integer range 0 to 3 :=2;
	variable timer_up_key : integer range 0 to 6 :=0;
	begin
		if RESET = '1' then
			Prescaler <= (others => '0');
			SquareX <= "1001010001";  
         SquareY <= "0110001011";
			flag_btn := '0';
			lock_key := 2;
			timer_up_key := 0;
		elsif rising_edge(CLK_24MHz) then
		   if (end_game = '0' and pause = '0') then
			Prescaler <= Prescaler + 1;	 
			if Prescaler = "0111010100110000000" then  
			if(Btn(0) = '0' or Btn(1) = '0') then  
			   flag_btn := '1';
				lock_key := 1;
					if(Btn(0) = '0') then flagR :='1'; flagL :='0';
					elsif(Btn(1) = '0') then flagL :='1'; flagR:='0'; 
					end if;				
			end if;
			
			
			if (lock_key = 1) then
			   timer_up_key := timer_up_key + 1;
			end if;
			
			if (timer_up_key = 5) then
			   timer_up_key := 0;
			   lock_key := 0;
		   end if;
			 
				if( lock_key = 1 )then
				   if(FlagR = '1') then
						if (SquareX - 2) > 110 then
							SquareX <= SquareX - 2;
					
						else
							Squarex <= Squarex;
						end if;
				   elsif(FlagL= '1') then
						if (SquareX + 2) < ((640-65)+21) then
							SquareX <= SquareX + 2;
					
						else
							Squarex<= Squarex;
						end if;
					else
				      SquareY <= SquareY;
			   	end if;	 
		   end if;		  
				Prescaler <= (others => '0');
			end if;
			end if;
		end if;
	end process square;		
	
shot: process(CLK_24MHz, RESET)
   variable flag_btn : bit:= '0';
	variable counter : integer := 1000;
	begin
		if RESET = '1' then
         flag_btn := '0';
			shotx <= SquareX + 6;
         shoty <= "0110001011";
		elsif rising_edge(CLK_24MHz) then
			if (end_game = '0' and pause = '0') then
				if (shoty <= 110) then 
				shotX <= SquareX + 6;
				shotY <= "0110001011";
				end if;
				if( Btn(0) = '0' or Btn(1) = '0')then
					 flag_btn := '1';
				end if;
				if(flag_btn = '1') then
					if( counter = 0 )then
						counter := 1000;
					end if;
					counter := counter - 1;
					
					if( counter = 0 )then  
						if(flag_btn = '1') then
							shotY <= shotY - 1;
						end if;	 
					end if;
				end if;
			end if;
		end if;
end process shot;
rock: process(CLK_24MHz, RESET)
   variable flag_btn,flagUP,FlagRight : bit:= '0';
	variable Z_Y,Z_x : integer range 0 to 6 := 3 ;
	variable counter : integer range 0 to 600001 :=600000;
	variable rand1 : integer range 0 to 5000 := 0;
	begin
	
		if RESET = '1' or rockflag = '0'  then
			rand1 := (random mod 5000) + 1;
			rockX <=std_logic_vector(to_unsigned(((rand1 mod 441) + 110),rockX'length));
         rockY <= "0001101110" ;
			Z_Y:= (rand1 mod 5) + 1;
			Z_X:= (5 - Z_X) + 1;
			counter := 600000;
			rocknum<= ((rand1/10) mod 5) + 4;
			if RESET = '1' then
			flag_btn := '0';	fast <= '0';	end if;
		elsif rising_edge(CLK_24MHz) then
		if (end_game = '0' and pause = '0') then
		if( Btn(0) = '0' or Btn(1) = '0')then
		    flag_btn := '1';
		end if;
		if( Btn(3) = '0')then
		    fast <= '1';
		end if;
		if(flag_btn = '1') then
			if( counter = 0 )then
				counter := 600000 - speed;
			end if;
		counter := counter - 1;			
			if( counter = 0 )then   
				if(flag_btn = '1') then
					if(rockx >= ((640-67)-21)) then flagUP :='1';
					elsif(rockx <= 111) then flagUp := '0';
					end if;
					if(rockY >= ((480-65)-21) ) then flagRight :='1';
					elsif(rocky <= 111) then flagright := '0';
					end if;
					if(flagUp='1') then rockX <= rockX - Z_X;
					elsif(flagUp='0') then rockX <= rockX + Z_X;
					end if;
					if(flagright='1') then rocky <= rocky - Z_y;
					elsif(flagright='0') then rocky <= rocky + Z_y;
					end if;
			   end if;	 

			end if;
		end if;
		end if;
		end if;
	end process rock;		
	process( CLK_24MHz, RESET)
	variable counter: integer:=9000000; 
	variable rock_num: integer range 0 to 9 := 0;
	variable flag: bit := '0';
	begin
	if RESET = '1' then
		lose <= '0';
		losegame <= '0';		
		score_signal <= 0;
		speed <= 100000 ;
		rock_num := 0;
	elsif( rising_edge(CLK_24MHz))then
		savedam <= rock_num;
		if(fast = '1') then
			speed <= 450000; end if;
		if ((SquareX > rockX AND SquareY > rocky AND SquareX < rockX+SquareWidth AND SquareY < rockY+SquareWidth) or 
		(SquareX+SquareWidth > rockX AND SquareY > rocky AND SquareX < rockX AND SquareY < rockY+SquareWidth)) then
			lose <= '1';
			loseGame <= '1';
		end if;
		if(flag = '1') then	counter := counter - 1 ; end if;
		if(counter = 0) then flag :='0'; end if;
		if (flag ='0' and(( shotX > rockX AND shotY > rocky AND shotx < rockX+SquareWidth AND shotY < rockY+SquareWidth) or
									(rockx > shotY and rockY > shotX and rockX <shotX+shotsize and rocky <shoty+shotsize ))) then
			rock_num := rock_num + 1;
			if(fast = '1') then
			score_signal <= score_signal + 4 ;
			else	score_signal <= score_signal + 1 ; end if;
			flag :='1';
			counter := 9000000;
			if(rocknum = rock_num) then
				rockflag <= '0';
				rock_num := 0;
				if(speed <= 450000) then
				speed <= speed + 100000; end if;
			end if;
				
			else rockflag <= '1';
			end if;
	end if;	
	end process;
	score <= score_signal;
	rockdam <= rocknum - savedam;
	rockmap <= rock8 when rockdam=8 
				else rock7 when rockdam=7
				else rock6 when rockdam=6
				else rock5 when rockdam=5
				else rock4 when rockdam=4
				else rock3 when rockdam=3
				else rock2 when rockdam=2
				else rock1 when rockdam=1
				else rock1;
	wall_color <= "101010" when end_game='0'
					else "110000" when losegame='1'
					else "001100";
   ColorOutput <= "110000" when losegame = '1' And end_game = '1' AND ScanlineX > 328 AND ScanlineY > 241 AND ScanlineX < 391 AND ScanlineY < 265 and endlose(CONV_INTEGER(scanlineY) mod 22 ,CONV_INTEGER (scanlinex) mod 66) = '1'
					else "001100" when losegame = '0' And end_game = '1' AND ScanlineX > 329 AND ScanlineY > 241 AND ScanlineX < 395 AND ScanlineY < 264 and endwin(CONV_INTEGER(scanlineY) mod 22 ,CONV_INTEGER (scanlinex) mod 66) = '1'
					else "111111" when  ScanlineX > rockX AND ScanlineY > rocky AND ScanlineX < rockX+SquareWidth AND ScanlineY < rockY+SquareWidth AND rockmap((CONV_INTEGER( scanlineY)-CONV_INTEGER(rockY)) mod 22 ,(CONV_INTEGER (scanlinex)-CONV_INTEGER(rockX)) mod 22) = '1'
					else  "111000" when  ScanlineX > rockX AND ScanlineY > rocky AND ScanlineX < rockX+SquareWidth AND ScanlineY < rockY+SquareWidth AND  rockmap ((CONV_INTEGER( scanlineY)-CONV_INTEGER(rockY)) mod 22 ,(CONV_INTEGER (scanlinex)-CONV_INTEGER(rockX)) mod 22) = '0'					
					else "010101" when ScanlineY < 480-62 AND ScanlineY > 480-87 And ScanlineX > ((640-65)+19) AND ScanlineX < ((640-65)+41) And home(CONV_INTEGER(scanlineY) mod 22 ,CONV_INTEGER (scanlinex) mod 22) = '1'
					else wall_color when ScanlineY < 480-62 AND ScanlineY > 480-87 And ScanlineX > ((640-65)+19) AND ScanlineX < ((640-65)+41) And home(CONV_INTEGER(scanlineY) mod 22 ,CONV_INTEGER (scanlinex) mod 22) = '0'
					else "011000" when  ScanlineX > SquareX AND ScanlineY > SquareY AND ScanlineX < SquareX+SquareWidth AND ScanlineY < SquareY+SquareWidth and tank((CONV_INTEGER( scanlineY)-CONV_INTEGER(SquareY)) mod 22 ,(CONV_INTEGER (scanlinex)-CONV_INTEGER(SquareX)) mod 22) = '1'
					else "000000" when  ScanlineX > SquareX AND ScanlineY > SquareY AND ScanlineX < SquareX+SquareWidth AND ScanlineY < SquareY+SquareWidth and tank((CONV_INTEGER( scanlineY)-CONV_INTEGER(SquareY)) mod 22 ,(CONV_INTEGER (scanlinex)-CONV_INTEGER(SquareX)) mod 22) = '0'		
					else "010101" when	ScanlineX > shotX AND ScanlineY > shoty AND ScanlineX < shotX+shotsize AND ScanlineY < shotY+Shotsize	AND shotmap((CONV_INTEGER( scanlineY)-CONV_INTEGER(shotY)) mod 22 ,(CONV_INTEGER (scanlinex)-CONV_INTEGER(shotX)) mod 7) = '1'
					else "000000" when 	ScanlineX > 110 AND ScanlineY > 110 AND ScanlineX < 640-68 AND ScanlineY < 480-62
					else "000000" when 	ScanlineY < 480-62 AND ScanlineY > 480-87 And ScanlineX >= 640-68 AND ScanlineX <= ((640-65)+19)
				   else "010101" when wall(CONV_INTEGER(scanlineY) mod 22 ,CONV_INTEGER (scanlinex) mod 22) = '1'
					else wall_color when wall(CONV_INTEGER(scanlineY) mod 22 ,CONV_INTEGER (scanlinex) mod 22) = '0'
					else	"000000" ;

	ColorOut <= ColorOutput;
end Behavioral;
